// ============================================================================
// Module: state_register
// Descrizione:
//   Questo modulo rappresenta un registro di stato parametrico per l'algoritmo 
//   ASCON (o simili), in grado di memorizzare e gestire 5 parole da 64 bit 
//   ciascuna (tipicamente lo stato interno dell'algoritmo).
//
//   Supporta due operazioni principali:
//     - **Scrittura parallela** dell'intero stato (`write_en`),
//     - **Shift seriale** dello stato, in due modalità:
//         • shift di PAR bit per parola (non mascherato),
//         • shift di (d+1)*PAR bit per parola (mascherato).
//
//   È progettato per integrarsi con architetture mascherate, adattandosi al 
//   grado di parallelismo e all’ordine di mascheramento specificato. Gestisce 
//   anche l’ultimo ciclo di shift con quantità inferiore di bit tramite `last_cycle`.
//
//   Parametri:
//     - COL_SIZE: numero di parole (default: 5),
//     - WORD_SIZE: dimensione in bit di ogni parola (default: 64),
//     - PAR: grado di parallelismo,
//     - d: ordine del mascheramento,
//     - SHIFT_PAR[_LAST], SHIFT_PAR_D_PLUS_1[_LAST]: gestiscono i casi di shift completi/parziali.
//
//   Output:
//     - `data_out`: stato completo attuale,
//     - `out_shifted_dplus1`: porzione di bit destinata allo shift mascherato.
//
// ============================================================================
import ascon_params::COL_SIZE;
import ascon_params::PAR;
import ascon_params::d;
import ascon_params::WORD_SIZE;
import ascon_params::SHIFT_PAR;
import ascon_params::SHIFT_PAR_D_PLUS_1;
import ascon_params::SHIFT_PAR_LAST;
import ascon_params::SHIFT_PAR_D_PLUS_1_LAST;

module state_register 
(
    input  logic clk,
    input  logic write_en,
    input  logic shift_en,
    input  logic shift_type, // 1 = shift 1, 0 = shift d+1
    input  logic last_cycle, 

    input  logic [COL_SIZE*WORD_SIZE-1:0] data_in,
    input  logic [COL_SIZE*SHIFT_PAR_D_PLUS_1-1:0] in_shifted_dplus1,
    input  logic [COL_SIZE*SHIFT_PAR-1:0]          in_shifted_1bit,
    
    output logic [COL_SIZE*SHIFT_PAR_D_PLUS_1-1:0] out_shifted_dplus1,
    output logic [COL_SIZE*WORD_SIZE-1:0] data_out
);

    logic [WORD_SIZE-1:0] state [0:COL_SIZE-1];
    (* keep = "true" *) logic [WORD_SIZE-1:0] next_state [0:COL_SIZE-1];

    generate 
    if (SHIFT_PAR_D_PLUS_1_LAST < WORD_SIZE) begin : gen_case1
        always_comb begin
            for (int i = 0; i < COL_SIZE; i++) begin
                next_state[i] = state[i]; // Default

                if (shift_en) begin
                    if (shift_type) begin
                        if (last_cycle) begin
                            // Ultimo ciclo con PAR_LAST
                            next_state[i] = {in_shifted_1bit[i*SHIFT_PAR +: SHIFT_PAR_LAST], state[i][WORD_SIZE-1:SHIFT_PAR_LAST]};
                        end else begin
                            // Cicli normali
                            next_state[i] = {in_shifted_1bit[i*SHIFT_PAR +: SHIFT_PAR], state[i][WORD_SIZE-1:SHIFT_PAR]};
                        end
                    end else begin
                        if (last_cycle) begin
                            next_state[i] = {in_shifted_dplus1[i*SHIFT_PAR_D_PLUS_1 +: SHIFT_PAR_D_PLUS_1_LAST], state[i][WORD_SIZE-1:SHIFT_PAR_D_PLUS_1_LAST]};
                        end else begin
                            next_state[i] = {in_shifted_dplus1[i*SHIFT_PAR_D_PLUS_1 +: SHIFT_PAR_D_PLUS_1], state[i][WORD_SIZE-1:SHIFT_PAR_D_PLUS_1]};
                        end
                    end
                end else if (write_en) begin
                    next_state[i] = data_in[i*WORD_SIZE +: WORD_SIZE];
                end
            end
        end

    end else begin : gen_case2
        always_comb begin
            for (int i = 0; i < COL_SIZE; i++) begin
                next_state[i] = state[i]; // Default

                if (shift_en) begin
                    if (shift_type) begin
                        if (last_cycle) begin
                            // Ultimo ciclo con PAR_LAST
                            next_state[i] = {in_shifted_1bit[i*SHIFT_PAR +: SHIFT_PAR_LAST], state[i][WORD_SIZE-1:SHIFT_PAR_LAST]};
                        end else begin
                            // Cicli normali
                            next_state[i] = {in_shifted_1bit[i*SHIFT_PAR +: SHIFT_PAR], state[i][WORD_SIZE-1:SHIFT_PAR]};
                        end
                    end else begin
                        // Ultimo ciclo con PAR_LAST
                        next_state[i] = in_shifted_dplus1[i*SHIFT_PAR_D_PLUS_1 +: WORD_SIZE];
                    end
                end else if (write_en) begin
                    next_state[i] = data_in[i*WORD_SIZE +: WORD_SIZE];
                end
            end
        end
    end
    endgenerate

    // === Blocco sequenziale
    always_ff @(posedge clk) begin
        for (int i = 0; i < COL_SIZE; i++) begin
            state[i] <= next_state[i];
        end
    end

    // === Output combinatorio
    generate
    if (SHIFT_PAR_D_PLUS_1_LAST < WORD_SIZE) begin : gen_caseNoPArMAx
        always_comb begin
            for (int i = 0; i < COL_SIZE; i++) begin
                out_shifted_dplus1[i*SHIFT_PAR_D_PLUS_1 +: SHIFT_PAR_D_PLUS_1] =
                state[i][SHIFT_PAR_D_PLUS_1-1:0];
                data_out[i*WORD_SIZE +: WORD_SIZE] = state[i];
            end
        end
    end
    else begin : gen_caseNoPArMAx
        always_comb begin
            for (int i = 0; i < COL_SIZE; i++) begin
                out_shifted_dplus1[i*WORD_SIZE +: WORD_SIZE] =
                state[i][WORD_SIZE-1:0];
                data_out[i*WORD_SIZE +: WORD_SIZE] = state[i];
            end
        end
    end
    endgenerate

endmodule
